module fewcore ();

endmodule

	